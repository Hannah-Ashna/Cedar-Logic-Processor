<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>383.433,-200.435,576.255,-297.537</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>418.5,-220</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_DECODER_2x4</type>
<position>431.5,-216.5</position>
<input>
<ID>ENABLE</ID>5 </input>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>40 </output>
<output>
<ID>OUT_2</ID>58 </output>
<output>
<ID>OUT_3</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_DECODER_2x4</type>
<position>431.5,-225</position>
<input>
<ID>ENABLE</ID>6 </input>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT_1</ID>20 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>EE_VDD</type>
<position>425.5,-215</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>EE_VDD</type>
<position>426.5,-223.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>DD_KEYPAD_HEX</type>
<position>419,-260.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>8 </output>
<output>
<ID>OUT_3</ID>7 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>438,-260.5</position>
<input>
<ID>ENABLE_0</ID>11 </input>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>7 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>14 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>443.5,-258</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>454,-259.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>464,-261</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>22</ID>
<type>DE_TO</type>
<position>472.5,-264.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>24</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>506,-257.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>16 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>472,-256.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>479,-258.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>488,-259.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>497,-260</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_REGISTER4</type>
<position>457,-233</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<input>
<ID>IN_2</ID>30 </input>
<input>
<ID>IN_3</ID>29 </input>
<output>
<ID>OUT_0</ID>24 </output>
<output>
<ID>OUT_1</ID>25 </output>
<output>
<ID>OUT_2</ID>26 </output>
<output>
<ID>OUT_3</ID>23 </output>
<input>
<ID>clear</ID>34 </input>
<input>
<ID>clock</ID>33 </input>
<input>
<ID>count_enable</ID>21 </input>
<input>
<ID>count_up</ID>22 </input>
<input>
<ID>load</ID>20 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>36</ID>
<type>FF_GND</type>
<position>457,-224</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>FF_GND</type>
<position>458,-225.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>463,-232.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>26 </input>
<input>
<ID>IN_3</ID>23 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>38 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>440,-234</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>443,-234.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>446,-235</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>448.5,-236</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>456,-242</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>48</ID>
<type>FF_GND</type>
<position>458,-238</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>475,-233.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>472.5,-234.5</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>470,-235.5</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>467,-236</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_REGISTER4</type>
<position>496,-233</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>48 </input>
<input>
<ID>IN_3</ID>47 </input>
<output>
<ID>OUT_0</ID>44 </output>
<output>
<ID>OUT_1</ID>45 </output>
<output>
<ID>OUT_2</ID>46 </output>
<output>
<ID>OUT_3</ID>43 </output>
<input>
<ID>clear</ID>52 </input>
<input>
<ID>clock</ID>51 </input>
<input>
<ID>count_enable</ID>41 </input>
<input>
<ID>count_up</ID>42 </input>
<input>
<ID>load</ID>57 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>57</ID>
<type>FF_GND</type>
<position>496,-224</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>FF_GND</type>
<position>497,-225.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>502,-232.5</position>
<input>
<ID>ENABLE_0</ID>58 </input>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>43 </input>
<output>
<ID>OUT_0</ID>56 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>54 </output>
<output>
<ID>OUT_3</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>479,-234</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>482,-234.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>485,-235</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>487.5,-236</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>495,-242</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>65</ID>
<type>FF_GND</type>
<position>497,-238</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_TO</type>
<position>514,-233.5</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>511.5,-234.5</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>68</ID>
<type>DE_TO</type>
<position>509,-235.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_TO</type>
<position>506,-236</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_REGISTER4</type>
<position>536,-233</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<input>
<ID>IN_2</ID>66 </input>
<input>
<ID>IN_3</ID>65 </input>
<output>
<ID>OUT_0</ID>62 </output>
<output>
<ID>OUT_1</ID>63 </output>
<output>
<ID>OUT_2</ID>64 </output>
<output>
<ID>OUT_3</ID>61 </output>
<input>
<ID>clear</ID>70 </input>
<input>
<ID>clock</ID>69 </input>
<input>
<ID>count_enable</ID>59 </input>
<input>
<ID>count_up</ID>60 </input>
<input>
<ID>load</ID>75 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>71</ID>
<type>FF_GND</type>
<position>536,-224</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>FF_GND</type>
<position>537,-225.5</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>542,-232.5</position>
<input>
<ID>ENABLE_0</ID>76 </input>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<input>
<ID>IN_2</ID>64 </input>
<input>
<ID>IN_3</ID>61 </input>
<output>
<ID>OUT_0</ID>74 </output>
<output>
<ID>OUT_1</ID>73 </output>
<output>
<ID>OUT_2</ID>72 </output>
<output>
<ID>OUT_3</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>519,-234</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>522,-234.5</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>525,-235</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>527.5,-236</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>535,-242</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>79</ID>
<type>FF_GND</type>
<position>537,-238</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>554,-233.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>551.5,-234.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>82</ID>
<type>DE_TO</type>
<position>549,-235.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>83</ID>
<type>DE_TO</type>
<position>546,-236</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>420,-242</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>424,-242</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423.5,-217,428.5,-217</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<connection>
<GID>4</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423.5,-218,428.5,-218</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>423.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>423.5,-219,423.5,-218</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>-218 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,-225.5,424.5,-221</points>
<intersection>-225.5 1</intersection>
<intersection>-221 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424.5,-225.5,428.5,-225.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423.5,-221,424.5,-221</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>424.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423.5,-226.5,428.5,-226.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>423.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>423.5,-226.5,423.5,-223</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>426.5,-215,428.5,-215</points>
<connection>
<GID>4</GID>
<name>ENABLE</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>427.5,-223.5,428.5,-223.5</points>
<connection>
<GID>6</GID>
<name>ENABLE</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436,-259,436,-257.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>424,-257.5,436,-257.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>436 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431,-260,436,-260</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>431 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>431,-260,431,-259.5</points>
<intersection>-260 1</intersection>
<intersection>-259.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>424,-259.5,431,-259.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>431 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431,-261,436,-261</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>431 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>431,-261.5,431,-261</points>
<intersection>-261.5 6</intersection>
<intersection>-261 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>424,-261.5,431,-261.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>431 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436,-263.5,436,-262</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-263.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>424,-263.5,436,-263.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>436 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438,-257.5,438,-218</points>
<connection>
<GID>14</GID>
<name>ENABLE_0</name></connection>
<intersection>-218 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-218,438,-218</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>438 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,-258,441.5,-258</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>440 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>440,-259,440,-258</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<intersection>-258 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,-259.5,452,-259.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>440 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>440,-260,440,-259.5</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<intersection>-259.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,-261,462,-261</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440,-264.5,440,-262</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>440,-264.5,470.5,-264.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>440 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474,-255.5,503,-255.5</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>474 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>474,-256.5,474,-255.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-255.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,-256.5,503,-256.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>481 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>481,-258.5,481,-256.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-256.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>490,-257.5,503,-257.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>490 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>490,-259.5,490,-257.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-257.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>499,-260,503,-260</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>503 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>503,-260,503,-258.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-260 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434.5,-225.5,456,-225.5</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>456 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>456,-228,456,-225.5</points>
<connection>
<GID>34</GID>
<name>load</name></connection>
<intersection>-225.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-228,457,-225</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<connection>
<GID>34</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,-228,458,-226.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<connection>
<GID>34</GID>
<name>count_up</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>461,-231,461,-231</points>
<connection>
<GID>34</GID>
<name>OUT_3</name></connection>
<connection>
<GID>40</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>461,-234,461,-234</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>461,-233,461,-233</points>
<connection>
<GID>34</GID>
<name>OUT_1</name></connection>
<connection>
<GID>40</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>461,-232,461,-232</points>
<connection>
<GID>34</GID>
<name>OUT_2</name></connection>
<connection>
<GID>40</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,-231,453,-231</points>
<connection>
<GID>34</GID>
<name>IN_3</name></connection>
<intersection>440 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>440,-232,440,-231</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-231 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>443,-232,453,-232</points>
<connection>
<GID>34</GID>
<name>IN_2</name></connection>
<intersection>443 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>443,-232.5,443,-232</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-232 1</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>446,-233,453,-233</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448.5,-234,453,-234</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-240,456,-237</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,-237,458,-237</points>
<connection>
<GID>34</GID>
<name>clear</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>475,-231.5,475,-231</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>465,-231,475,-231</points>
<connection>
<GID>40</GID>
<name>OUT_3</name></connection>
<intersection>475 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>472.5,-232.5,472.5,-232</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-232 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>465,-232,472.5,-232</points>
<connection>
<GID>40</GID>
<name>OUT_2</name></connection>
<intersection>472.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-233.5,470,-233</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-233 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>465,-233,470,-233</points>
<connection>
<GID>40</GID>
<name>OUT_1</name></connection>
<intersection>470 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>465,-234,467,-234</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,-229.5,463,-217</points>
<connection>
<GID>40</GID>
<name>ENABLE_0</name></connection>
<intersection>-217 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-217,463,-217</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>463 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496,-228,496,-225</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-228,497,-226.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>count_up</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>500,-231,500,-231</points>
<connection>
<GID>56</GID>
<name>OUT_3</name></connection>
<connection>
<GID>59</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>500,-234,500,-234</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>500,-233,500,-233</points>
<connection>
<GID>56</GID>
<name>OUT_1</name></connection>
<connection>
<GID>59</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>500,-232,500,-232</points>
<connection>
<GID>56</GID>
<name>OUT_2</name></connection>
<connection>
<GID>59</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>479,-231,492,-231</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>479 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>479,-232,479,-231</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-231 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>482,-232,492,-232</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>482 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>482,-232.5,482,-232</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-232 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>485,-233,492,-233</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>487.5,-234,492,-234</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495,-240,495,-237</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-237,497,-237</points>
<connection>
<GID>56</GID>
<name>clear</name></connection>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-231.5,514,-231</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>504,-231,514,-231</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-232.5,511.5,-232</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-232 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>504,-232,511.5,-232</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,-233.5,509,-233</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-233 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>504,-233,509,-233</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>509 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>504,-234,506,-234</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495,-228,495,-224.5</points>
<connection>
<GID>56</GID>
<name>load</name></connection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-224.5,495,-224.5</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>495 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,-229.5,502,-216</points>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<intersection>-216 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-216,502,-216</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>536,-228,536,-225</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<connection>
<GID>70</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,-228,537,-226.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<connection>
<GID>70</GID>
<name>count_up</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,-231,540,-231</points>
<connection>
<GID>70</GID>
<name>OUT_3</name></connection>
<connection>
<GID>73</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,-234,540,-234</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,-233,540,-233</points>
<connection>
<GID>70</GID>
<name>OUT_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,-232,540,-232</points>
<connection>
<GID>70</GID>
<name>OUT_2</name></connection>
<connection>
<GID>73</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-231,532,-231</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>519 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>519,-232,519,-231</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-231 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,-232,532,-232</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>522 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>522,-232.5,522,-232</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-232 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>525,-233,532,-233</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527.5,-234,532,-234</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535,-240,535,-237</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>537,-237,537,-237</points>
<connection>
<GID>70</GID>
<name>clear</name></connection>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>554,-231.5,554,-231</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>544,-231,554,-231</points>
<connection>
<GID>73</GID>
<name>OUT_3</name></connection>
<intersection>554 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>551.5,-232.5,551.5,-232</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>-232 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>544,-232,551.5,-232</points>
<connection>
<GID>73</GID>
<name>OUT_2</name></connection>
<intersection>551.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>549,-233.5,549,-233</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-233 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>544,-233,549,-233</points>
<connection>
<GID>73</GID>
<name>OUT_1</name></connection>
<intersection>549 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>544,-234,546,-234</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434.5,-223.5,535,-223.5</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>535 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535,-228,535,-223.5</points>
<connection>
<GID>70</GID>
<name>load</name></connection>
<intersection>-223.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542,-229.5,542,-215</points>
<connection>
<GID>73</GID>
<name>ENABLE_0</name></connection>
<intersection>-215 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-215,542,-215</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>542 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422,-242,422,-242</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>502.371,-5.56966,1896.37,-707.57</PageViewport></page 1>
<page 2>
<PageViewport>-16.1536,657.815,1377.85,-44.1852</PageViewport></page 2>
<page 3>
<PageViewport>5.99978,659.231,1400,-42.7693</PageViewport></page 3>
<page 4>
<PageViewport>285.701,7.53383,1679.7,-694.466</PageViewport></page 4>
<page 5>
<PageViewport>110.435,85.1829,1504.44,-616.817</PageViewport></page 5>
<page 6>
<PageViewport>-657.666,883.549,736.334,181.549</PageViewport></page 6>
<page 7>
<PageViewport>-0.000223028,659.231,1394,-42.7693</PageViewport></page 7>
<page 8>
<PageViewport>-0.000223028,659.231,1394,-42.7693</PageViewport></page 8>
<page 9>
<PageViewport>-0.000223028,659.231,1394,-42.7693</PageViewport></page 9></circuit>