<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-2156.37,566.913,-2069.94,523.39</PageViewport>
<gate>
<ID>1</ID>
<type>BA_NAND2</type>
<position>-2126,547</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>-2126,540</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_NAND2</type>
<position>-2104,547</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>-2104,540</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>-2093,547</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>-2093,540</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-2150,551</position>
<gparam>LABEL_TEXT Data</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-2150,540</position>
<gparam>LABEL_TEXT Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>-2093,549</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-2093,542</position>
<gparam>LABEL_TEXT Not Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>BA_NAND2</type>
<position>-2114,548</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>-2114,539</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-2121.5,555.5</position>
<gparam>LABEL_TEXT Master Slave Circuit - NAND Gates</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>-2135,548</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND2</type>
<position>-2135,539</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>-2150,549</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>-2121,551.5</position>
<input>
<ID>N_in2</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>-2150,538</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2143,534</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>-2121,535.5</position>
<input>
<ID>N_in3</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2141,540</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2111,548,-2107,548</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2111,539,-2107,539</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>4</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2097,540,-2097,544</points>
<intersection>540 2</intersection>
<intersection>544 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2107,544,-2097,544</points>
<intersection>-2107 3</intersection>
<intersection>-2097 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2101,540,-2094,540</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-2097 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2107,544,-2107,546</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>544 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2096,543,-2096,547</points>
<intersection>543 2</intersection>
<intersection>547 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2101,547,-2094,547</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>-2096 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2107,543,-2096,543</points>
<intersection>-2107 3</intersection>
<intersection>-2096 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2107,541,-2107,543</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>543 2</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2120,538,-2120,544</points>
<intersection>538 5</intersection>
<intersection>540 2</intersection>
<intersection>544 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2129,544,-2120,544</points>
<intersection>-2129 3</intersection>
<intersection>-2120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2123,540,-2120,540</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-2120 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2129,544,-2129,546</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>544 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-2121,538,-2117,538</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-2121 6</intersection>
<intersection>-2120 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-2121,536.5,-2121,538</points>
<connection>
<GID>22</GID>
<name>N_in3</name></connection>
<intersection>538 5</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2121,543,-2121,550.5</points>
<connection>
<GID>18</GID>
<name>N_in2</name></connection>
<intersection>543 2</intersection>
<intersection>547 1</intersection>
<intersection>549 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2123,547,-2121,547</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>-2121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2129,543,-2121,543</points>
<intersection>-2129 3</intersection>
<intersection>-2121 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2129,541,-2129,543</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>543 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-2121,549,-2117,549</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-2121 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2148,549,-2138,549</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-2146 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-2146,540,-2146,549</points>
<intersection>540 8</intersection>
<intersection>549 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-2146,540,-2143,540</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-2146 7</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2148,538,-2138,538</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-2145 4</intersection>
<intersection>-2144 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-2144,538,-2144,547</points>
<intersection>538 1</intersection>
<intersection>547 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2144,547,-2138,547</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-2144 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-2145,534,-2145,538</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>538 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2132,548,-2129,548</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2132,539,-2129,539</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2118,534,-2118,547</points>
<intersection>534 2</intersection>
<intersection>540 3</intersection>
<intersection>547 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2141,534,-2118,534</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-2118 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-2118,540,-2117,540</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-2118 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-2118,547,-2117,547</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-2118 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2139,540,-2138,540</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>50.4894,-26.478,127.311,-65.1642</PageViewport></page 1>
<page 2>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>-2.14686,3.46927e-006,179.947,-91.7</PageViewport></page 9></circuit>