<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-2146.93,561.478,-2083.64,528.837</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-2126,550</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-2126,541</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>-2114,549</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>-2114,542</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>-2103,549</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>-2103,542</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-2126,552</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>-2126,543</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-2103,551</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-2103,544</position>
<gparam>LABEL_TEXT Not Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-2113,555.5</position>
<gparam>LABEL_TEXT S-R Latch - NAND Gates</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2124,550,-2117,550</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-2117 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-2117,550,-2117,550</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>550 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2124,541,-2117,541</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-2117 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-2117,541,-2117,541</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>541 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2107,542,-2107,546</points>
<intersection>542 2</intersection>
<intersection>542 2</intersection>
<intersection>546 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2117,546,-2107,546</points>
<intersection>-2117 3</intersection>
<intersection>-2107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2111,542,-2104,542</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>-2107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2117,546,-2117,548</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>546 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2106,545,-2106,549</points>
<intersection>545 2</intersection>
<intersection>549 1</intersection>
<intersection>549 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2111,549,-2104,549</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>-2106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2117,545,-2106,545</points>
<intersection>-2117 3</intersection>
<intersection>-2106 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2117,543,-2117,545</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>545 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>51.3953,-26.4781,126.405,-65.1641</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 9></circuit>