<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-2149.83,561.478,-2085.02,528.837</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-2140,551</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-2140,540</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_NAND2</type>
<position>-2115,549</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>-2115,542</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>-2104,549</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>-2104,542</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-2140,553.5</position>
<gparam>LABEL_TEXT Data</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-2140,542.5</position>
<gparam>LABEL_TEXT Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>-2104,551</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-2104,544</position>
<gparam>LABEL_TEXT Not Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>-2131,550</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>-2131,541</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-2121,557</position>
<gparam>LABEL_TEXT D-Latch with Enable - NAND Gates</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2128,550,-2118,550</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-2125 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-2125,546,-2125,550</points>
<intersection>546 3</intersection>
<intersection>550 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2134,546,-2125,546</points>
<intersection>-2134 4</intersection>
<intersection>-2125 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-2134,542,-2134,546</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>546 3</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2128,541,-2118,541</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2108,542,-2108,546</points>
<intersection>542 2</intersection>
<intersection>546 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2118,546,-2108,546</points>
<intersection>-2118 3</intersection>
<intersection>-2108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2112,542,-2105,542</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-2108 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2118,546,-2118,548</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>546 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2107,545,-2107,549</points>
<intersection>545 2</intersection>
<intersection>549 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2112,549,-2105,549</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>-2107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2118,545,-2107,545</points>
<intersection>-2118 3</intersection>
<intersection>-2107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2118,543,-2118,545</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>545 2</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2138,540,-2134,540</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-2136 2</intersection>
<intersection>-2134 7</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-2136,540,-2136,549</points>
<intersection>540 1</intersection>
<intersection>549 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2136,549,-2134,549</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-2136 2</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-2134,540,-2134,540</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>540 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2138,551,-2134,551</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-2134 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-2134,551,-2134,551</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>551 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>50.4895,-26.478,127.311,-65.1642</PageViewport></page 1>
<page 2>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>-2.14686,2.31285e-006,179.947,-91.7</PageViewport></page 9></circuit>