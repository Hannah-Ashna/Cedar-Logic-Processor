<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-31.942,9.03254,145.347,-80.248</PageViewport>
<gate>
<ID>1</ID>
<type>BA_DECODER_2x4</type>
<position>43,-33.5</position>
<input>
<ID>ENABLE</ID>85 </input>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT_0</ID>76 </output>
<output>
<ID>OUT_1</ID>14 </output>
<output>
<ID>OUT_2</ID>52 </output>
<output>
<ID>OUT_3</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_REGISTER4</type>
<position>25,-29.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>54 </input>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>59 </output>
<output>
<ID>OUT_3</ID>58 </output>
<input>
<ID>clear</ID>16 </input>
<input>
<ID>clock</ID>53 </input>
<input>
<ID>count_enable</ID>15 </input>
<input>
<ID>count_up</ID>15 </input>
<input>
<ID>load</ID>67 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_DECODER_2x4</type>
<position>44,-27</position>
<input>
<ID>ENABLE</ID>85 </input>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT_0</ID>17 </output>
<output>
<ID>OUT_1</ID>18 </output>
<output>
<ID>OUT_2</ID>51 </output>
<output>
<ID>OUT_3</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>52,-65</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>61,-66</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>70.5,-67</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>79,-68</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>71,-63</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>81,-64</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>90.5,-65</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>100,-66</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>82,-49</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>79.5,-49</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>77,-49</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>84.5,-49</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>56,-50</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>58,-50</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>60.5,-50</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>62.5,-50</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_REGISTER4</type>
<position>102.5,-44</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>48 </input>
<input>
<ID>IN_3</ID>47 </input>
<output>
<ID>OUT_0</ID>41 </output>
<output>
<ID>OUT_1</ID>39 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>38 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>42 </input>
<input>
<ID>count_enable</ID>36 </input>
<input>
<ID>count_up</ID>35 </input>
<input>
<ID>load</ID>52 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>21</ID>
<type>FF_GND</type>
<position>103.5,-38</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>FF_GND</type>
<position>102.5,-36.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>FF_GND</type>
<position>103.5,-49</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>109,-43.5</position>
<input>
<ID>ENABLE_0</ID>51 </input>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>38 </input>
<output>
<ID>OUT_0</ID>43 </output>
<output>
<ID>OUT_1</ID>44 </output>
<output>
<ID>OUT_2</ID>45 </output>
<output>
<ID>OUT_3</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>101.5,-50</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>117,-47</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>114.5,-47</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>112,-47</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>119.5,-47</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>91,-48</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>93,-48</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>95.5,-48</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>97.5,-48</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>88.5,-6.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>109,-14</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>109,-11.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>109,-9</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>109,-17</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>39</ID>
<type>FF_GND</type>
<position>25,-21.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>FF_GND</type>
<position>26,-35.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>24,-42.5</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>42</ID>
<type>DD_KEYPAD_HEX</type>
<position>35,-66</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>106.5,-65</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>23 </input>
<input>
<ID>IN_3</ID>24 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>44</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>47.5,-66.5</position>
<input>
<ID>ENABLE_0</ID>17 </input>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>22 </output>
<output>
<ID>OUT_1</ID>21 </output>
<output>
<ID>OUT_2</ID>20 </output>
<output>
<ID>OUT_3</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_REGISTER4</type>
<position>67.5,-46</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>33 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>31 </input>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>10 </output>
<output>
<ID>OUT_3</ID>8 </output>
<input>
<ID>clear</ID>7 </input>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>count_enable</ID>6 </input>
<input>
<ID>count_up</ID>5 </input>
<input>
<ID>load</ID>14 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>46</ID>
<type>FF_GND</type>
<position>68.5,-40</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>FF_GND</type>
<position>67.5,-38.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>FF_GND</type>
<position>68.5,-51</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>74,-45.5</position>
<input>
<ID>ENABLE_0</ID>18 </input>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT_0</ID>27 </output>
<output>
<ID>OUT_1</ID>28 </output>
<output>
<ID>OUT_2</ID>29 </output>
<output>
<ID>OUT_3</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>66.5,-52.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>24.5,3.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>7,-39</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>9,-39</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>11.5,-39</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>13.5,-39</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>14,-16.5</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AE_DFF_LOW</type>
<position>11.5,-10.5</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUTINV_0</ID>62 </output>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clear</ID>66 </input>
<input>
<ID>clock</ID>63 </input>
<input>
<ID>set</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>59</ID>
<type>DA_FROM</type>
<position>3.5,-11.5</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>60</ID>
<type>DE_TO</type>
<position>18,-8.5</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>61</ID>
<type>EE_VDD</type>
<position>11.5,-5.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>EE_VDD</type>
<position>11.5,-15.5</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>11,-23</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_REGISTER4</type>
<position>89.5,-22</position>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>70 </output>
<output>
<ID>OUT_2</ID>69 </output>
<output>
<ID>OUT_3</ID>68 </output>
<input>
<ID>clear</ID>73 </input>
<input>
<ID>clock</ID>72 </input>
<input>
<ID>count_enable</ID>75 </input>
<input>
<ID>count_up</ID>74 </input>
<input>
<ID>load</ID>88 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_RAM_4x4</type>
<position>99.5,-11.5</position>
<input>
<ID>ADDRESS_0</ID>71 </input>
<input>
<ID>ADDRESS_1</ID>70 </input>
<input>
<ID>ADDRESS_2</ID>69 </input>
<input>
<ID>ADDRESS_3</ID>68 </input>
<input>
<ID>DATA_IN_0</ID>80 </input>
<input>
<ID>DATA_IN_1</ID>81 </input>
<input>
<ID>DATA_IN_2</ID>82 </input>
<input>
<ID>DATA_IN_3</ID>83 </input>
<output>
<ID>DATA_OUT_0</ID>80 </output>
<output>
<ID>DATA_OUT_1</ID>81 </output>
<output>
<ID>DATA_OUT_2</ID>82 </output>
<output>
<ID>DATA_OUT_3</ID>83 </output>
<input>
<ID>ENABLE_0</ID>86 </input>
<input>
<ID>write_clock</ID>78 </input>
<input>
<ID>write_enable</ID>79 </input>
<gparam>angle 90</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 1</lparam>
<lparam>Address:1 6</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>88.5,-28</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>67</ID>
<type>FF_GND</type>
<position>90.5,-27</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>EE_VDD</type>
<position>90.5,-14.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>85,-12.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>42.5,3.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_SMALL_INVERTER</type>
<position>47,3.5</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>53.5,3.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>37.5,-21</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_OR2</type>
<position>60.5,-4</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BB_CLOCK</type>
<position>18.5,3.5</position>
<output>
<ID>CLK</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>93.5,-27</position>
<gparam>LABEL_TEXT Program counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>49.5,-38</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>80,-17</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-63,45.5,-63</points>
<connection>
<GID>42</GID>
<name>OUT_3</name></connection>
<intersection>45.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45.5,-65,45.5,-63</points>
<connection>
<GID>44</GID>
<name>IN_3</name></connection>
<intersection>-63 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-66,40.5,-65</points>
<intersection>-66 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-66,45.5,-66</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-65,40.5,-65</points>
<connection>
<GID>42</GID>
<name>OUT_2</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-67,45.5,-67</points>
<connection>
<GID>42</GID>
<name>OUT_1</name></connection>
<intersection>45.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>45.5,-67,45.5,-67</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-69,40.5,-68</points>
<intersection>-69 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-68,45.5,-68</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-69,40.5,-69</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>68.5,-41,68.5,-41</points>
<connection>
<GID>45</GID>
<name>count_up</name></connection>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-41,67.5,-39.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<connection>
<GID>45</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>68.5,-50,68.5,-50</points>
<connection>
<GID>45</GID>
<name>clear</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71.5,-44,72,-44</points>
<connection>
<GID>49</GID>
<name>IN_3</name></connection>
<connection>
<GID>45</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71.5,-46,72,-46</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<connection>
<GID>45</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71.5,-45,72,-45</points>
<connection>
<GID>49</GID>
<name>IN_2</name></connection>
<connection>
<GID>45</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71.5,-47,72,-47</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>66.5,-50.5,66.5,-50</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,3.5,22.5,3.5</points>
<connection>
<GID>76</GID>
<name>CLK</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-41,66.5,-34</points>
<connection>
<GID>45</GID>
<name>load</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-34,66.5,-34</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-24.5,25,-22.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>count_enable</name></connection>
<intersection>-24.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>25,-24.5,26,-24.5</points>
<connection>
<GID>2</GID>
<name>count_up</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>26,-34.5,26,-33.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-63.5,47.5,-28.5</points>
<connection>
<GID>44</GID>
<name>ENABLE_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-28.5,47.5,-28.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-42.5,74,-27.5</points>
<connection>
<GID>49</GID>
<name>ENABLE_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-27.5,74,-27.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>49.5,-65,50,-65</points>
<connection>
<GID>44</GID>
<name>OUT_3</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-66,59,-66</points>
<connection>
<GID>44</GID>
<name>OUT_2</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-67,68.5,-67</points>
<connection>
<GID>44</GID>
<name>OUT_1</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-68,77,-68</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-64,103.5,-64</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-63,103.5,-63</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92.5,-65,103.5,-65</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102,-66,103.5,-66</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-47,77,-47</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-47,79.5,-46</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-46,79.5,-46</points>
<connection>
<GID>49</GID>
<name>OUT_1</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-47,82,-45</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-45,82,-45</points>
<connection>
<GID>49</GID>
<name>OUT_2</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-47,84.5,-44</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-44,84.5,-44</points>
<connection>
<GID>49</GID>
<name>OUT_3</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-48,56,-44</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-44,63.5,-44</points>
<connection>
<GID>45</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-48,58,-45</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-45,63.5,-45</points>
<connection>
<GID>45</GID>
<name>IN_2</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-48,60.5,-46</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-46,63.5,-46</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-48,62.5,-47</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-47,63.5,-47</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-39,103.5,-39</points>
<connection>
<GID>20</GID>
<name>count_up</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-39,102.5,-37.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>103.5,-48,103.5,-48</points>
<connection>
<GID>20</GID>
<name>clear</name></connection>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>106.5,-42,107,-42</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<connection>
<GID>20</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>106.5,-44,107,-44</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>106.5,-43,107,-43</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<connection>
<GID>20</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>106.5,-45,107,-45</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>101.5,-48,101.5,-48</points>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-45,112,-45</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-45,114.5,-44</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-44,114.5,-44</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-45,117,-43</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-43,117,-43</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-45,119.5,-42</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-42,119.5,-42</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-46,91,-42</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-42,98.5,-42</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-46,93,-43</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-43,98.5,-43</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-46,95.5,-44</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-44,98.5,-44</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-46,97.5,-45</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-45,98.5,-45</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-40.5,109,-34</points>
<connection>
<GID>24</GID>
<name>ENABLE_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-34,109,-34</points>
<intersection>76.5 2</intersection>
<intersection>109 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76.5,-34,76.5,-26.5</points>
<intersection>-34 1</intersection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-26.5,76.5,-26.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>76.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-39,75,-33</points>
<intersection>-39 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-33,75,-33</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-39,101.5,-39</points>
<connection>
<GID>20</GID>
<name>load</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>24,-40.5,24,-33.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-37,7,-27.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-27.5,21,-27.5</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-37,9,-28.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-28.5,21,-28.5</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-37,11.5,-29.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-29.5,21,-29.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-37,13.5,-30.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-30.5,21,-30.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-27.5,41,-27.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-28.5,41,-28.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-35,35.5,-30.5</points>
<intersection>-35 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-30.5,35.5,-30.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-35,40,-35</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-34,36.5,-29.5</points>
<intersection>-34 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-29.5,36.5,-29.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-34,40,-34</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-11.5,26.5,-1.5</points>
<intersection>-11.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-11.5,26.5,-11.5</points>
<connection>
<GID>58</GID>
<name>OUTINV_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-1.5,26.5,-1.5</points>
<intersection>3 3</intersection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>3,-8.5,3,-1.5</points>
<intersection>-8.5 4</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>3,-8.5,8.5,-8.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>3 3</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-11.5,8.5,-11.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<connection>
<GID>58</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-8.5,16,-8.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-6.5,11.5,-6.5</points>
<connection>
<GID>58</GID>
<name>set</name></connection>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-14.5,11.5,-14.5</points>
<connection>
<GID>58</GID>
<name>clear</name></connection>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-24.5,24,-23</points>
<connection>
<GID>2</GID>
<name>load</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-23,24,-23</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-20,98,-16.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_3</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-20,98,-20</points>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-21,99,-16.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_2</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-21,99,-21</points>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-22,100,-16.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_1</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-22,100,-22</points>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-23,101,-16.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-23,101,-23</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-26,88.5,-26</points>
<connection>
<GID>64</GID>
<name>clock</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-26,90.5,-26</points>
<connection>
<GID>64</GID>
<name>clear</name></connection>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-17,90.5,-15.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<connection>
<GID>64</GID>
<name>count_up</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-17,89.5,-12.5</points>
<connection>
<GID>64</GID>
<name>count_enable</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-12.5,89.5,-12.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-38,46,-35</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-38,47.5,-38</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,3.5,45,3.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>45 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>45,-3,45,3.5</points>
<intersection>-3 9</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>45,-3,57.5,-3</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>45 8</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-6.5,98,-6.5</points>
<connection>
<GID>65</GID>
<name>write_clock</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-6.5,99,-5</points>
<connection>
<GID>65</GID>
<name>write_enable</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-5,99,-5</points>
<intersection>70 2</intersection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>70,-32,70,-5</points>
<intersection>-32 3</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>46,-32,70,-32</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>70 2</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-10,104.5,-9</points>
<connection>
<GID>65</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>65</GID>
<name>DATA_IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-9,107,-9</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11.5,104.5,-11</points>
<connection>
<GID>65</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>65</GID>
<name>DATA_IN_1</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-11.5,107,-11.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-14,105.5,-12</points>
<intersection>-14 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-14,107,-14</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-12,105.5,-12</points>
<connection>
<GID>65</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>65</GID>
<name>DATA_IN_2</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-17,104.5,-13</points>
<connection>
<GID>65</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>65</GID>
<name>DATA_IN_3</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-17,107,-17</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,3.5,51.5,3.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-32,40,-21</points>
<connection>
<GID>1</GID>
<name>ENABLE</name></connection>
<intersection>-25.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-21,40,-21</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-25.5,41,-25.5</points>
<connection>
<GID>3</GID>
<name>ENABLE</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63.5,-4,100,-4</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>100 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>100,-6.5,100,-4</points>
<connection>
<GID>65</GID>
<name>ENABLE_0</name></connection>
<intersection>-4 1</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-25.5,52,-5</points>
<intersection>-25.5 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-5,57.5,-5</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-25.5,52,-25.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-17,88.5,-17</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>88.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>88.5,-17,88.5,-17</points>
<connection>
<GID>64</GID>
<name>load</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 1>
<page 2>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 2>
<page 3>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 3>
<page 4>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 4>
<page 5>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 5>
<page 6>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 6>
<page 7>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 7>
<page 8>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 8>
<page 9>
<PageViewport>0,92.302,996.133,-409.337</PageViewport></page 9></circuit>